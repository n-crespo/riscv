`timescale 1ns / 1ps
// Decodes 32-bit RISC-V instructions into standard fields
module decoder (
    input  [31:0] instr,
    output [ 6:0] opcode,
    output [ 4:0] rd,
    output [ 2:0] funct3,
    output [ 4:0] rs1,
    output [ 4:0] rs2,
    output [ 6:0] funct7
);

  // slice the instruction into its respective components based on RISC-V architecture
  assign opcode = instr[6:0];
  assign rd     = instr[11:7];
  assign funct3 = instr[14:12];
  assign rs1    = instr[19:15];
  assign rs2    = instr[24:20];
  assign funct7 = instr[31:25];

endmodule
